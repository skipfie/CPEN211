module tb_task1(output err);
  // your implementation here
endmodule: tb_task1
