module tb_idecoder(output err);
  // your implementation here
endmodule: tb_idecoder
