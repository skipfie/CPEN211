module task2(input clk, input rst_n, input [7:0] start_pc, output[15:0] out);
    // how to do ldr
    /*
    ldr 1:
    reg_sel = 10
    en_A = 1

    ldr 2:
    sel_A = 0
    sel_B = 1
    en_C = 1
    
    ldr 3:
    load_addr = 1

    ldr 4:
    sel_addr = 0

    ldr 5:
    wb_sel = 11
    reg_sel = 01
    w_en = 1


    */
endmodule: task2
