module tb_cpu(output err);
  // your implementation here
endmodule: tb_cpu
