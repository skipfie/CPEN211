module task1(input clk, input rst_n, input [7:0] start_pc, output[15:0] out);
  // your implementation here
endmodule: task1
