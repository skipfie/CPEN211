module tb_shifter(output err);
    reg shift_in 
endmodule: tb_shifter
