module task2(input clk, input rst_n, input [7:0] start_pc, output[15:0] out);
    // how to do ldr
    /*
    ldr 1:
    

    */
endmodule: task2
