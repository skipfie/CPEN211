module tb_datapath(output err);
  reg 


  initial begin
    

    $stop;
  end

endmodule: tb_datapath
