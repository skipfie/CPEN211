module tb_controller(output err);
  // your implementation here
endmodule: tb_controller
